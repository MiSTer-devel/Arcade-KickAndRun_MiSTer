
localparam CORE_CLK_SYS = 72;
localparam CORE_CLK_6 = (CORE_CLK_SYS/6)-1;
localparam CORE_CLK_4 = (CORE_CLK_SYS/4)-1;
localparam CORE_CLK_1 = (CORE_CLK_SYS/1)-1;
